
`timescale 1fs/1fs
module ctle_tb;

    real vdd;
    real vss;
    real vinp;
    real voutp;
    real vinn;
    real voutn;
    integer get_value_file_file;

    

    ctle #(
        
    ) dut (
        .vdd(vdd),
        .vss(vss),
        .vinp(vinp),
        .voutp(voutp),
        .vinn(vinn),
        .voutn(voutn)
    );

    initial begin
        get_value_file_file = $fopen("/home/dstanley/research/fixture_demo/build/get_value_file.txt", "w");
        vdd <= 1.8;
        #(0*1s);
        vss <= 0;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8859382209404254;
        #(0*1s);
        vinn <= 0.9207223413512122;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9152890571351513;
        #(0*1s);
        vinn <= 0.8913715051564863;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9112893869874528;
        #(0*1s);
        vinn <= 0.9157220098663337;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.936405450941883;
        #(0*1s);
        vinn <= 0.8906059459119035;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8983947265591615;
        #(0*1s);
        vinn <= 0.9427077324765732;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9365015596928463;
        #(0*1s);
        vinn <= 0.9046008993428885;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8854665655433138;
        #(0*1s);
        vinn <= 0.9322551233783813;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9329152153350821;
        #(0*1s);
        vinn <= 0.884806473586613;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9135356913669516;
        #(0*1s);
        vinn <= 0.9466167395209636;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9454022113735691;
        #(0*1s);
        vinn <= 0.9147502195143461;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9195031604342003;
        #(0*1s);
        vinn <= 0.9330625837550124;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9465332205559288;
        #(0*1s);
        vinn <= 0.9060325236332839;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9234715570944307;
        #(0*1s);
        vinn <= 0.9714835301210138;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9671087782295958;
        #(0*1s);
        vinn <= 0.9278463089858487;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9217958338138267;
        #(0*1s);
        vinn <= 0.9685179244137704;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9685616961926206;
        #(0*1s);
        vinn <= 0.9217520620349765;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9219413609306275;
        #(0*1s);
        vinn <= 0.9588420497567278;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9567778029055556;
        #(0*1s);
        vinn <= 0.9240056077817997;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8933397804873966;
        #(0*1s);
        vinn <= 0.9221573681206567;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9234890874502335;
        #(0*1s);
        vinn <= 0.8920080611578198;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.906901072032982;
        #(0*1s);
        vinn <= 0.9527152173145736;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9489066341569966;
        #(0*1s);
        vinn <= 0.910709655190559;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9009372343678432;
        #(0*1s);
        vinn <= 0.9459251122694354;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9380129186956297;
        #(0*1s);
        vinn <= 0.9088494279416489;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8928112170203896;
        #(0*1s);
        vinn <= 0.9422554627010974;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9424379175781705;
        #(0*1s);
        vinn <= 0.8926287621433164;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.894944574576996;
        #(0*1s);
        vinn <= 0.9367065875380162;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9318559827075847;
        #(0*1s);
        vinn <= 0.8997951794074275;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9269231081217383;
        #(0*1s);
        vinn <= 0.9515288899218423;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9620637756887805;
        #(0*1s);
        vinn <= 0.9163882223548;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9313836253119102;
        #(0*1s);
        vinn <= 0.9371493936774561;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9575275635826831;
        #(0*1s);
        vinn <= 0.9110054554066832;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9293120321718616;
        #(0*1s);
        vinn <= 0.9681759204538148;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9706624730292346;
        #(0*1s);
        vinn <= 0.9268254795964419;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8964685874395859;
        #(0*1s);
        vinn <= 0.9432761648752286;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9291228400311056;
        #(0*1s);
        vinn <= 0.9106219122837089;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8760141674347892;
        #(0*1s);
        vinn <= 0.9240662325411049;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9248439413830467;
        #(0*1s);
        vinn <= 0.8752364585928474;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9229961814223785;
        #(0*1s);
        vinn <= 0.961637681555317;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9634914225105081;
        #(0*1s);
        vinn <= 0.9211424404671874;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9240902445162678;
        #(0*1s);
        vinn <= 0.9437836490721077;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9527418005870063;
        #(0*1s);
        vinn <= 0.9151320930013691;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9013067560203311;
        #(0*1s);
        vinn <= 0.9500182954858384;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9412345778032162;
        #(0*1s);
        vinn <= 0.9100904737029533;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.9128276249739152;
        #(0*1s);
        vinn <= 0.9619867329690569;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9460579935787665;
        #(0*1s);
        vinn <= 0.9287563643642056;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8922369592256489;
        #(0*1s);
        vinn <= 0.9313591119521571;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9366376192634162;
        #(0*1s);
        vinn <= 0.8869584519143899;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", vinn);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1e-09*1s);
        vinp <= 0.8805631716320353;
        #(0*1s);
        vinn <= 0.9274895616179654;
        #(0*1s);
        #(1e-09*1s);
        vinp <= 0.9261033694325713;
        #(0*1s);
        vinn <= 0.8819493638174294;
        #(0*1s);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutp);
        $fwrite(get_value_file_file, "%0.15f\n", $realtime/1s);//\n", voutn);
        #(1.1000000000000001e-09*1s);
        $fclose(get_value_file_file);

        #20 $finish;
    end

endmodule
